module stack_mem();
