module sign_extension (
