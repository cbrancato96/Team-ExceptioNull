module cpu()
  
  wire [7:0] pc
